//--------------------------------------------------------------------------
//  Data memory test bench
//--------------------------------------------------------------------------

module datamemorytest();
    reg clk, address, writeEnable, dataIn;
    wire dataOut;

