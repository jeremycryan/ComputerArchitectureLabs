`define AND and #30
`define XOR xor #50
//Instruction Fetch Unit which outputs an address
//to Instruction Memory and is able to jump and
//branch when provided appropriate control signals

module ifu
(
    output[29:0] address,
    output[31:0] pcStore,
    input[25:0] targetInstr,
    input[15:0] imm16,
    input[31:0] jRrs,
    input branch,jump, zero, bne, jl, jr, clk
);

reg[31:0] pc;
wire[31:0] immExtend;
wire[31:0] addend;
wire[31:0] sum;
wire[31:0] concatenate;
wire[31:0] pcNext;
wire[31:0] addendInter;
wire[31:0] jumpAddress;

wire do_branch, branch_condition;

initial begin
    pc <= 32'b00000000000000000000000000000000;
end

assign pcStore = sum;

assign address = pc[29:0];
signExtend1632 extend(immExtend,imm16);
`XOR condition(branch_condition,zero,bne); // Takes care of BNE and BEQ
`AND branchy(do_branch,branch,branch_condition); // Decides if to branch
mux2_32 addMux1(addendInter,32'b00000000000000000000000000000000,immExtend,do_branch);
mux2_32 addMux2(addend,addendInter,32'b1,jl);
Adder32Bit adder(
    .sum(sum),
    .carryout(),
    .a(pc),
    .b(addend),
    .carryin(1'b1)
);

assign concatenate = {pc[31:28],targetInstr};
mux2_32 jumpMux1(jumpAddress, concatenate, jRrs, jr);
mux2_32 jumpMux2(pcNext,jumpAddress,sum,jump); 

// Assign pc to pcNext on clk edge
always @(posedge clk)begin
    pc <= pcNext;
end

endmodule
