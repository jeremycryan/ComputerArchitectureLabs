//  full lst

`define AND and #50
`define OR or #50
`define NOT not #50

module FullSLT(
    output out,
    input a,
    input b,
    input prev
);
