`include "sign_extend.v"

module signExtend1632Test();
    
    // Stuff here

endmodule
